module decoder4to16
  (
	input [3:0] w, 
	input En,         
	output reg [15:0] y  
  );

	always @(*) begin
		case ({En, w})  
			5'b10000: y = 16'b0000000000000001;
			5'b10001: y = 16'b0000000000000010;
			5'b10010: y = 16'b0000000000000100;
			5'b10011: y = 16'b0000000000001000;
			5'b10100: y = 16'b0000000000010000;
			5'b10101: y = 16'b0000000000100000;
			5'b10110: y = 16'b0000000001000000;
			5'b10111: y = 16'b0000000010000000;
			5'b11000: y = 16'b0000000100000000;
			default:  y = 16'b0000000000000000;  
		endcase
	end

endmodule
